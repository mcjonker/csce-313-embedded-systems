// nios_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,       //       clk.clk
		input  wire        reset_reset_n, //     reset.reset_n
		output wire [12:0] sdram_addr,    //     sdram.addr
		output wire [1:0]  sdram_ba,      //          .ba
		output wire        sdram_cas_n,   //          .cas_n
		output wire        sdram_cke,     //          .cke
		output wire        sdram_cs_n,    //          .cs_n
		inout  wire [31:0] sdram_dq,      //          .dq
		output wire [3:0]  sdram_dqm,     //          .dqm
		output wire        sdram_ras_n,   //          .ras_n
		output wire        sdram_we_n,    //          .we_n
		output wire        sdram_clk_clk, // sdram_clk.clk
		inout  wire [15:0] sram_DQ,       //      sram.DQ
		output wire [19:0] sram_ADDR,     //          .ADDR
		output wire        sram_LB_N,     //          .LB_N
		output wire        sram_UB_N,     //          .UB_N
		output wire        sram_CE_N,     //          .CE_N
		output wire        sram_OE_N,     //          .OE_N
		output wire        sram_WE_N,     //          .WE_N
		output wire        vga_CLK,       //       vga.CLK
		output wire        vga_HS,        //          .HS
		output wire        vga_VS,        //          .VS
		output wire        vga_BLANK,     //          .BLANK
		output wire        vga_SYNC,      //          .SYNC
		output wire [7:0]  vga_R,         //          .R
		output wire [7:0]  vga_G,         //          .G
		output wire [7:0]  vga_B          //          .B
	);

	wire         video_alpha_blender_0_avalon_blended_source_valid;                                        // video_alpha_blender_0:output_valid -> dual_clock_fifo:stream_in_valid
	wire  [29:0] video_alpha_blender_0_avalon_blended_source_data;                                         // video_alpha_blender_0:output_data -> dual_clock_fifo:stream_in_data
	wire         video_alpha_blender_0_avalon_blended_source_ready;                                        // dual_clock_fifo:stream_in_ready -> video_alpha_blender_0:output_ready
	wire         video_alpha_blender_0_avalon_blended_source_startofpacket;                                // video_alpha_blender_0:output_startofpacket -> dual_clock_fifo:stream_in_startofpacket
	wire         video_alpha_blender_0_avalon_blended_source_endofpacket;                                  // video_alpha_blender_0:output_endofpacket -> dual_clock_fifo:stream_in_endofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_valid;                               // video_character_buffer_with_dma_0:stream_valid -> video_alpha_blender_0:foreground_valid
	wire  [39:0] video_character_buffer_with_dma_0_avalon_char_source_data;                                // video_character_buffer_with_dma_0:stream_data -> video_alpha_blender_0:foreground_data
	wire         video_character_buffer_with_dma_0_avalon_char_source_ready;                               // video_alpha_blender_0:foreground_ready -> video_character_buffer_with_dma_0:stream_ready
	wire         video_character_buffer_with_dma_0_avalon_char_source_startofpacket;                       // video_character_buffer_with_dma_0:stream_startofpacket -> video_alpha_blender_0:foreground_startofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_endofpacket;                         // video_character_buffer_with_dma_0:stream_endofpacket -> video_alpha_blender_0:foreground_endofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_valid;                                            // dual_clock_fifo:stream_out_valid -> vga:valid
	wire  [29:0] dual_clock_fifo_avalon_dc_buffer_source_data;                                             // dual_clock_fifo:stream_out_data -> vga:data
	wire         dual_clock_fifo_avalon_dc_buffer_source_ready;                                            // vga:ready -> dual_clock_fifo:stream_out_ready
	wire         dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                                    // dual_clock_fifo:stream_out_startofpacket -> vga:startofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                                      // dual_clock_fifo:stream_out_endofpacket -> vga:endofpacket
	wire         dma_buffer_avalon_pixel_source_valid;                                                     // dma_buffer:stream_valid -> rgb_resampler:stream_in_valid
	wire  [23:0] dma_buffer_avalon_pixel_source_data;                                                      // dma_buffer:stream_data -> rgb_resampler:stream_in_data
	wire         dma_buffer_avalon_pixel_source_ready;                                                     // rgb_resampler:stream_in_ready -> dma_buffer:stream_ready
	wire         dma_buffer_avalon_pixel_source_startofpacket;                                             // dma_buffer:stream_startofpacket -> rgb_resampler:stream_in_startofpacket
	wire         dma_buffer_avalon_pixel_source_endofpacket;                                               // dma_buffer:stream_endofpacket -> rgb_resampler:stream_in_endofpacket
	wire         rgb_resampler_avalon_rgb_source_valid;                                                    // rgb_resampler:stream_out_valid -> video_scaler:stream_in_valid
	wire  [29:0] rgb_resampler_avalon_rgb_source_data;                                                     // rgb_resampler:stream_out_data -> video_scaler:stream_in_data
	wire         rgb_resampler_avalon_rgb_source_ready;                                                    // video_scaler:stream_in_ready -> rgb_resampler:stream_out_ready
	wire         rgb_resampler_avalon_rgb_source_startofpacket;                                            // rgb_resampler:stream_out_startofpacket -> video_scaler:stream_in_startofpacket
	wire         rgb_resampler_avalon_rgb_source_endofpacket;                                              // rgb_resampler:stream_out_endofpacket -> video_scaler:stream_in_endofpacket
	wire         sys_sdram_pll_sys_clk_clk;                                                                // sys_sdram_pll:sys_clk_clk -> [avalon_st_adapter:in_clk_0_clk, dma_buffer:clk, dual_clock_fifo:clk_stream_in, irq_mapper:clk, jtag:clk, mm_interconnect_0:sys_sdram_pll_sys_clk_clk, processor:clk, rgb_resampler:clk, rst_controller_001:clk, rst_controller_002:clk, rst_controller_004:clk, rst_controller_005:clk, sram_controller:clk, sysid_qsys_0:clock, timer_0:clk, video_alpha_blender_0:clk, video_character_buffer_with_dma_0:clk, video_scaler:clk]
	wire         video_pll_0_vga_clk_clk;                                                                  // video_pll_0:vga_clk_clk -> [dual_clock_fifo:clk_stream_out, rst_controller_003:clk, rst_controller_008:clk, vga:clk]
	wire         processor_custom_instruction_master_readra;                                               // processor:E_ci_combo_readra -> processor_custom_instruction_master_translator:ci_slave_readra
	wire         processor_custom_instruction_master_readrb;                                               // processor:E_ci_combo_readrb -> processor_custom_instruction_master_translator:ci_slave_readrb
	wire   [4:0] processor_custom_instruction_master_multi_b;                                              // processor:A_ci_multi_b -> processor_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] processor_custom_instruction_master_multi_c;                                              // processor:A_ci_multi_c -> processor_custom_instruction_master_translator:ci_slave_multi_c
	wire         processor_custom_instruction_master_reset_req;                                            // processor:A_ci_multi_reset_req -> processor_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] processor_custom_instruction_master_multi_a;                                              // processor:A_ci_multi_a -> processor_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] processor_custom_instruction_master_result;                                               // processor_custom_instruction_master_translator:ci_slave_result -> processor:E_ci_combo_result
	wire  [31:0] processor_custom_instruction_master_datab;                                                // processor:E_ci_combo_datab -> processor_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] processor_custom_instruction_master_dataa;                                                // processor:E_ci_combo_dataa -> processor_custom_instruction_master_translator:ci_slave_dataa
	wire         processor_custom_instruction_master_writerc;                                              // processor:E_ci_combo_writerc -> processor_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] processor_custom_instruction_master_multi_dataa;                                          // processor:A_ci_multi_dataa -> processor_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         processor_custom_instruction_master_multi_writerc;                                        // processor:A_ci_multi_writerc -> processor_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [4:0] processor_custom_instruction_master_a;                                                    // processor:E_ci_combo_a -> processor_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] processor_custom_instruction_master_b;                                                    // processor:E_ci_combo_b -> processor_custom_instruction_master_translator:ci_slave_b
	wire  [31:0] processor_custom_instruction_master_multi_result;                                         // processor_custom_instruction_master_translator:ci_slave_multi_result -> processor:A_ci_multi_result
	wire         processor_custom_instruction_master_clk;                                                  // processor:A_ci_multi_clock -> processor_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] processor_custom_instruction_master_multi_datab;                                          // processor:A_ci_multi_datab -> processor_custom_instruction_master_translator:ci_slave_multi_datab
	wire   [4:0] processor_custom_instruction_master_c;                                                    // processor:E_ci_combo_c -> processor_custom_instruction_master_translator:ci_slave_c
	wire  [31:0] processor_custom_instruction_master_ipending;                                             // processor:E_ci_combo_ipending -> processor_custom_instruction_master_translator:ci_slave_ipending
	wire         processor_custom_instruction_master_start;                                                // processor:A_ci_multi_start -> processor_custom_instruction_master_translator:ci_slave_multi_start
	wire         processor_custom_instruction_master_done;                                                 // processor_custom_instruction_master_translator:ci_slave_multi_done -> processor:A_ci_multi_done
	wire   [7:0] processor_custom_instruction_master_n;                                                    // processor:E_ci_combo_n -> processor_custom_instruction_master_translator:ci_slave_n
	wire         processor_custom_instruction_master_estatus;                                              // processor:E_ci_combo_estatus -> processor_custom_instruction_master_translator:ci_slave_estatus
	wire         processor_custom_instruction_master_clk_en;                                               // processor:A_ci_multi_clk_en -> processor_custom_instruction_master_translator:ci_slave_multi_clken
	wire         processor_custom_instruction_master_reset;                                                // processor:A_ci_multi_reset -> processor_custom_instruction_master_translator:ci_slave_multi_reset
	wire         processor_custom_instruction_master_multi_readrb;                                         // processor:A_ci_multi_readrb -> processor_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         processor_custom_instruction_master_multi_readra;                                         // processor:A_ci_multi_readra -> processor_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] processor_custom_instruction_master_multi_n;                                              // processor:A_ci_multi_n -> processor_custom_instruction_master_translator:ci_slave_multi_n
	wire  [31:0] processor_custom_instruction_master_translator_comb_ci_master_result;                     // processor_custom_instruction_master_comb_xconnect:ci_slave_result -> processor_custom_instruction_master_translator:comb_ci_master_result
	wire         processor_custom_instruction_master_translator_comb_ci_master_readra;                     // processor_custom_instruction_master_translator:comb_ci_master_readra -> processor_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] processor_custom_instruction_master_translator_comb_ci_master_a;                          // processor_custom_instruction_master_translator:comb_ci_master_a -> processor_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] processor_custom_instruction_master_translator_comb_ci_master_b;                          // processor_custom_instruction_master_translator:comb_ci_master_b -> processor_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         processor_custom_instruction_master_translator_comb_ci_master_readrb;                     // processor_custom_instruction_master_translator:comb_ci_master_readrb -> processor_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] processor_custom_instruction_master_translator_comb_ci_master_c;                          // processor_custom_instruction_master_translator:comb_ci_master_c -> processor_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         processor_custom_instruction_master_translator_comb_ci_master_estatus;                    // processor_custom_instruction_master_translator:comb_ci_master_estatus -> processor_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] processor_custom_instruction_master_translator_comb_ci_master_ipending;                   // processor_custom_instruction_master_translator:comb_ci_master_ipending -> processor_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] processor_custom_instruction_master_translator_comb_ci_master_datab;                      // processor_custom_instruction_master_translator:comb_ci_master_datab -> processor_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] processor_custom_instruction_master_translator_comb_ci_master_dataa;                      // processor_custom_instruction_master_translator:comb_ci_master_dataa -> processor_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         processor_custom_instruction_master_translator_comb_ci_master_writerc;                    // processor_custom_instruction_master_translator:comb_ci_master_writerc -> processor_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] processor_custom_instruction_master_translator_comb_ci_master_n;                          // processor_custom_instruction_master_translator:comb_ci_master_n -> processor_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] processor_custom_instruction_master_comb_xconnect_ci_master0_result;                      // processor_custom_instruction_master_comb_slave_translator0:ci_slave_result -> processor_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         processor_custom_instruction_master_comb_xconnect_ci_master0_readra;                      // processor_custom_instruction_master_comb_xconnect:ci_master0_readra -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] processor_custom_instruction_master_comb_xconnect_ci_master0_a;                           // processor_custom_instruction_master_comb_xconnect:ci_master0_a -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] processor_custom_instruction_master_comb_xconnect_ci_master0_b;                           // processor_custom_instruction_master_comb_xconnect:ci_master0_b -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         processor_custom_instruction_master_comb_xconnect_ci_master0_readrb;                      // processor_custom_instruction_master_comb_xconnect:ci_master0_readrb -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] processor_custom_instruction_master_comb_xconnect_ci_master0_c;                           // processor_custom_instruction_master_comb_xconnect:ci_master0_c -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         processor_custom_instruction_master_comb_xconnect_ci_master0_estatus;                     // processor_custom_instruction_master_comb_xconnect:ci_master0_estatus -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] processor_custom_instruction_master_comb_xconnect_ci_master0_ipending;                    // processor_custom_instruction_master_comb_xconnect:ci_master0_ipending -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] processor_custom_instruction_master_comb_xconnect_ci_master0_datab;                       // processor_custom_instruction_master_comb_xconnect:ci_master0_datab -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] processor_custom_instruction_master_comb_xconnect_ci_master0_dataa;                       // processor_custom_instruction_master_comb_xconnect:ci_master0_dataa -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         processor_custom_instruction_master_comb_xconnect_ci_master0_writerc;                     // processor_custom_instruction_master_comb_xconnect:ci_master0_writerc -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] processor_custom_instruction_master_comb_xconnect_ci_master0_n;                           // processor_custom_instruction_master_comb_xconnect:ci_master0_n -> processor_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] processor_custom_instruction_master_comb_slave_translator0_ci_master_result;              // nios_custom_instr_floating_point_2_0:s1_result -> processor_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] processor_custom_instruction_master_comb_slave_translator0_ci_master_datab;               // processor_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s1_datab
	wire  [31:0] processor_custom_instruction_master_comb_slave_translator0_ci_master_dataa;               // processor_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s1_dataa
	wire   [3:0] processor_custom_instruction_master_comb_slave_translator0_ci_master_n;                   // processor_custom_instruction_master_comb_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s1_n
	wire         processor_custom_instruction_master_translator_multi_ci_master_readra;                    // processor_custom_instruction_master_translator:multi_ci_master_readra -> processor_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] processor_custom_instruction_master_translator_multi_ci_master_a;                         // processor_custom_instruction_master_translator:multi_ci_master_a -> processor_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] processor_custom_instruction_master_translator_multi_ci_master_b;                         // processor_custom_instruction_master_translator:multi_ci_master_b -> processor_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         processor_custom_instruction_master_translator_multi_ci_master_clk;                       // processor_custom_instruction_master_translator:multi_ci_master_clk -> processor_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         processor_custom_instruction_master_translator_multi_ci_master_readrb;                    // processor_custom_instruction_master_translator:multi_ci_master_readrb -> processor_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] processor_custom_instruction_master_translator_multi_ci_master_c;                         // processor_custom_instruction_master_translator:multi_ci_master_c -> processor_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         processor_custom_instruction_master_translator_multi_ci_master_start;                     // processor_custom_instruction_master_translator:multi_ci_master_start -> processor_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         processor_custom_instruction_master_translator_multi_ci_master_reset_req;                 // processor_custom_instruction_master_translator:multi_ci_master_reset_req -> processor_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         processor_custom_instruction_master_translator_multi_ci_master_done;                      // processor_custom_instruction_master_multi_xconnect:ci_slave_done -> processor_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] processor_custom_instruction_master_translator_multi_ci_master_n;                         // processor_custom_instruction_master_translator:multi_ci_master_n -> processor_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] processor_custom_instruction_master_translator_multi_ci_master_result;                    // processor_custom_instruction_master_multi_xconnect:ci_slave_result -> processor_custom_instruction_master_translator:multi_ci_master_result
	wire         processor_custom_instruction_master_translator_multi_ci_master_clk_en;                    // processor_custom_instruction_master_translator:multi_ci_master_clken -> processor_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] processor_custom_instruction_master_translator_multi_ci_master_datab;                     // processor_custom_instruction_master_translator:multi_ci_master_datab -> processor_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] processor_custom_instruction_master_translator_multi_ci_master_dataa;                     // processor_custom_instruction_master_translator:multi_ci_master_dataa -> processor_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         processor_custom_instruction_master_translator_multi_ci_master_reset;                     // processor_custom_instruction_master_translator:multi_ci_master_reset -> processor_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         processor_custom_instruction_master_translator_multi_ci_master_writerc;                   // processor_custom_instruction_master_translator:multi_ci_master_writerc -> processor_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_readra;                     // processor_custom_instruction_master_multi_xconnect:ci_master0_readra -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master0_a;                          // processor_custom_instruction_master_multi_xconnect:ci_master0_a -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master0_b;                          // processor_custom_instruction_master_multi_xconnect:ci_master0_b -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_readrb;                     // processor_custom_instruction_master_multi_xconnect:ci_master0_readrb -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master0_c;                          // processor_custom_instruction_master_multi_xconnect:ci_master0_c -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_clk;                        // processor_custom_instruction_master_multi_xconnect:ci_master0_clk -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_ipending;                   // processor_custom_instruction_master_multi_xconnect:ci_master0_ipending -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_start;                      // processor_custom_instruction_master_multi_xconnect:ci_master0_start -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_reset_req;                  // processor_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_done;                       // processor_custom_instruction_master_multi_slave_translator0:ci_slave_done -> processor_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] processor_custom_instruction_master_multi_xconnect_ci_master0_n;                          // processor_custom_instruction_master_multi_xconnect:ci_master0_n -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_result;                     // processor_custom_instruction_master_multi_slave_translator0:ci_slave_result -> processor_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_estatus;                    // processor_custom_instruction_master_multi_xconnect:ci_master0_estatus -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                     // processor_custom_instruction_master_multi_xconnect:ci_master0_clken -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_datab;                      // processor_custom_instruction_master_multi_xconnect:ci_master0_datab -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_dataa;                      // processor_custom_instruction_master_multi_xconnect:ci_master0_dataa -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_reset;                      // processor_custom_instruction_master_multi_xconnect:ci_master0_reset -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_writerc;                    // processor_custom_instruction_master_multi_xconnect:ci_master0_writerc -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator0_ci_master_result;             // nios_custom_instr_floating_point_2_0:s2_result -> processor_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_clk;                // processor_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_2_0:s2_clk
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;             // processor_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_2_0:s2_clk_en
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator0_ci_master_datab;              // processor_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s2_datab
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator0_ci_master_dataa;              // processor_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s2_dataa
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_start;              // processor_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_2_0:s2_start
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_reset;              // processor_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_2_0:s2_reset
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_reset_req;          // processor_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios_custom_instr_floating_point_2_0:s2_reset_req
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_done;               // nios_custom_instr_floating_point_2_0:s2_done -> processor_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] processor_custom_instruction_master_multi_slave_translator0_ci_master_n;                  // processor_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s2_n
	wire         dma_buffer_avalon_pixel_dma_master_waitrequest;                                           // mm_interconnect_0:dma_buffer_avalon_pixel_dma_master_waitrequest -> dma_buffer:master_waitrequest
	wire  [31:0] dma_buffer_avalon_pixel_dma_master_readdata;                                              // mm_interconnect_0:dma_buffer_avalon_pixel_dma_master_readdata -> dma_buffer:master_readdata
	wire  [31:0] dma_buffer_avalon_pixel_dma_master_address;                                               // dma_buffer:master_address -> mm_interconnect_0:dma_buffer_avalon_pixel_dma_master_address
	wire         dma_buffer_avalon_pixel_dma_master_read;                                                  // dma_buffer:master_read -> mm_interconnect_0:dma_buffer_avalon_pixel_dma_master_read
	wire         dma_buffer_avalon_pixel_dma_master_readdatavalid;                                         // mm_interconnect_0:dma_buffer_avalon_pixel_dma_master_readdatavalid -> dma_buffer:master_readdatavalid
	wire         dma_buffer_avalon_pixel_dma_master_lock;                                                  // dma_buffer:master_arbiterlock -> mm_interconnect_0:dma_buffer_avalon_pixel_dma_master_lock
	wire  [31:0] processor_data_master_readdata;                                                           // mm_interconnect_0:processor_data_master_readdata -> processor:d_readdata
	wire         processor_data_master_waitrequest;                                                        // mm_interconnect_0:processor_data_master_waitrequest -> processor:d_waitrequest
	wire         processor_data_master_debugaccess;                                                        // processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:processor_data_master_debugaccess
	wire  [28:0] processor_data_master_address;                                                            // processor:d_address -> mm_interconnect_0:processor_data_master_address
	wire   [3:0] processor_data_master_byteenable;                                                         // processor:d_byteenable -> mm_interconnect_0:processor_data_master_byteenable
	wire         processor_data_master_read;                                                               // processor:d_read -> mm_interconnect_0:processor_data_master_read
	wire         processor_data_master_readdatavalid;                                                      // mm_interconnect_0:processor_data_master_readdatavalid -> processor:d_readdatavalid
	wire         processor_data_master_write;                                                              // processor:d_write -> mm_interconnect_0:processor_data_master_write
	wire  [31:0] processor_data_master_writedata;                                                          // processor:d_writedata -> mm_interconnect_0:processor_data_master_writedata
	wire  [31:0] processor_instruction_master_readdata;                                                    // mm_interconnect_0:processor_instruction_master_readdata -> processor:i_readdata
	wire         processor_instruction_master_waitrequest;                                                 // mm_interconnect_0:processor_instruction_master_waitrequest -> processor:i_waitrequest
	wire  [28:0] processor_instruction_master_address;                                                     // processor:i_address -> mm_interconnect_0:processor_instruction_master_address
	wire         processor_instruction_master_read;                                                        // processor:i_read -> mm_interconnect_0:processor_instruction_master_read
	wire         processor_instruction_master_readdatavalid;                                               // mm_interconnect_0:processor_instruction_master_readdatavalid -> processor:i_readdatavalid
	wire  [15:0] mm_interconnect_0_sram_controller_avalon_sram_slave_readdata;                             // sram_controller:readdata -> mm_interconnect_0:sram_controller_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_controller_avalon_sram_slave_address;                              // mm_interconnect_0:sram_controller_avalon_sram_slave_address -> sram_controller:address
	wire         mm_interconnect_0_sram_controller_avalon_sram_slave_read;                                 // mm_interconnect_0:sram_controller_avalon_sram_slave_read -> sram_controller:read
	wire   [1:0] mm_interconnect_0_sram_controller_avalon_sram_slave_byteenable;                           // mm_interconnect_0:sram_controller_avalon_sram_slave_byteenable -> sram_controller:byteenable
	wire         mm_interconnect_0_sram_controller_avalon_sram_slave_readdatavalid;                        // sram_controller:readdatavalid -> mm_interconnect_0:sram_controller_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_controller_avalon_sram_slave_write;                                // mm_interconnect_0:sram_controller_avalon_sram_slave_write -> sram_controller:write
	wire  [15:0] mm_interconnect_0_sram_controller_avalon_sram_slave_writedata;                            // mm_interconnect_0:sram_controller_avalon_sram_slave_writedata -> sram_controller:writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata;    // video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest; // video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address;     // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read;        // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata;   // video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address;    // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	wire   [3:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write;      // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	wire  [31:0] mm_interconnect_0_dma_buffer_avalon_control_slave_readdata;                               // dma_buffer:slave_readdata -> mm_interconnect_0:dma_buffer_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_dma_buffer_avalon_control_slave_address;                                // mm_interconnect_0:dma_buffer_avalon_control_slave_address -> dma_buffer:slave_address
	wire         mm_interconnect_0_dma_buffer_avalon_control_slave_read;                                   // mm_interconnect_0:dma_buffer_avalon_control_slave_read -> dma_buffer:slave_read
	wire   [3:0] mm_interconnect_0_dma_buffer_avalon_control_slave_byteenable;                             // mm_interconnect_0:dma_buffer_avalon_control_slave_byteenable -> dma_buffer:slave_byteenable
	wire         mm_interconnect_0_dma_buffer_avalon_control_slave_write;                                  // mm_interconnect_0:dma_buffer_avalon_control_slave_write -> dma_buffer:slave_write
	wire  [31:0] mm_interconnect_0_dma_buffer_avalon_control_slave_writedata;                              // mm_interconnect_0:dma_buffer_avalon_control_slave_writedata -> dma_buffer:slave_writedata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                                      // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                                        // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                                     // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                                         // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                                            // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                                           // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                                       // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_rgb_resampler_avalon_rgb_slave_readdata;                                // rgb_resampler:slave_readdata -> mm_interconnect_0:rgb_resampler_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_rgb_resampler_avalon_rgb_slave_read;                                    // mm_interconnect_0:rgb_resampler_avalon_rgb_slave_read -> rgb_resampler:slave_read
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                                    // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                                     // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_processor_debug_mem_slave_readdata;                                     // processor:debug_mem_slave_readdata -> mm_interconnect_0:processor_debug_mem_slave_readdata
	wire         mm_interconnect_0_processor_debug_mem_slave_waitrequest;                                  // processor:debug_mem_slave_waitrequest -> mm_interconnect_0:processor_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_processor_debug_mem_slave_debugaccess;                                  // mm_interconnect_0:processor_debug_mem_slave_debugaccess -> processor:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_processor_debug_mem_slave_address;                                      // mm_interconnect_0:processor_debug_mem_slave_address -> processor:debug_mem_slave_address
	wire         mm_interconnect_0_processor_debug_mem_slave_read;                                         // mm_interconnect_0:processor_debug_mem_slave_read -> processor:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_processor_debug_mem_slave_byteenable;                                   // mm_interconnect_0:processor_debug_mem_slave_byteenable -> processor:debug_mem_slave_byteenable
	wire         mm_interconnect_0_processor_debug_mem_slave_write;                                        // mm_interconnect_0:processor_debug_mem_slave_write -> processor:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_processor_debug_mem_slave_writedata;                                    // mm_interconnect_0:processor_debug_mem_slave_writedata -> processor:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;                                         // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;                                           // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;                                        // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;                                            // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                                               // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;                                         // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;                                      // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;                                              // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;                                          // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                                  // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                                    // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                                     // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                                       // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                                   // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                                                                 // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                 // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] processor_irq_irq;                                                                        // irq_mapper:sender_irq -> processor:irq
	wire         video_scaler_avalon_scaler_source_valid;                                                  // video_scaler:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] video_scaler_avalon_scaler_source_data;                                                   // video_scaler:stream_out_data -> avalon_st_adapter:in_0_data
	wire         video_scaler_avalon_scaler_source_ready;                                                  // avalon_st_adapter:in_0_ready -> video_scaler:stream_out_ready
	wire   [1:0] video_scaler_avalon_scaler_source_channel;                                                // video_scaler:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         video_scaler_avalon_scaler_source_startofpacket;                                          // video_scaler:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         video_scaler_avalon_scaler_source_endofpacket;                                            // video_scaler:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                                            // avalon_st_adapter:out_0_valid -> video_alpha_blender_0:background_valid
	wire  [29:0] avalon_st_adapter_out_0_data;                                                             // avalon_st_adapter:out_0_data -> video_alpha_blender_0:background_data
	wire         avalon_st_adapter_out_0_ready;                                                            // video_alpha_blender_0:background_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                                                    // avalon_st_adapter:out_0_startofpacket -> video_alpha_blender_0:background_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                                      // avalon_st_adapter:out_0_endofpacket -> video_alpha_blender_0:background_endofpacket
	wire         rst_controller_reset_out_reset;                                                           // rst_controller:reset_out -> [rst_controller_004:reset_in0, rst_controller_008:reset_in0]
	wire         sys_sdram_pll_reset_source_reset;                                                         // sys_sdram_pll:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in2, rst_controller_005:reset_in2, rst_controller_006:reset_in1, rst_controller_007:reset_in1, rst_controller_008:reset_in2]
	wire         rst_controller_001_reset_out_reset;                                                       // rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, dma_buffer:reset, mm_interconnect_0:dma_buffer_reset_reset_bridge_in_reset_reset, rgb_resampler:reset, sram_controller:reset, video_alpha_blender_0:reset, video_character_buffer_with_dma_0:reset, video_scaler:reset]
	wire         rst_controller_002_reset_out_reset;                                                       // rst_controller_002:reset_out -> dual_clock_fifo:reset_stream_in
	wire         video_pll_0_reset_source_reset;                                                           // video_pll_0:reset_source_reset -> rst_controller_002:reset_in0
	wire         rst_controller_003_reset_out_reset;                                                       // rst_controller_003:reset_out -> dual_clock_fifo:reset_stream_out
	wire         rst_controller_004_reset_out_reset;                                                       // rst_controller_004:reset_out -> [jtag:rst_n, mm_interconnect_0:jtag_reset_reset_bridge_in_reset_reset, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire         rst_controller_005_reset_out_reset;                                                       // rst_controller_005:reset_out -> [irq_mapper:reset, mm_interconnect_0:processor_reset_reset_bridge_in_reset_reset, processor:reset_n]
	wire         rst_controller_005_reset_out_reset_req;                                                   // rst_controller_005:reset_req -> [processor:reset_req, rst_translator:reset_req_in]
	wire         processor_debug_reset_request_reset;                                                      // processor:debug_reset_request -> rst_controller_005:reset_in1
	wire         rst_controller_006_reset_out_reset;                                                       // rst_controller_006:reset_out -> [mm_interconnect_0:sdram_controller_reset_reset_bridge_in_reset_reset, sdram_controller:reset_n]
	wire         rst_controller_007_reset_out_reset;                                                       // rst_controller_007:reset_out -> [sys_sdram_pll:ref_reset_reset, video_pll_0:ref_reset_reset]
	wire         rst_controller_008_reset_out_reset;                                                       // rst_controller_008:reset_out -> vga:reset

	nios_system_dma_buffer dma_buffer (
		.clk                  (sys_sdram_pll_sys_clk_clk),                                    //                     clk.clk
		.reset                (rst_controller_001_reset_out_reset),                           //                   reset.reset
		.master_readdatavalid (dma_buffer_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (dma_buffer_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (dma_buffer_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (dma_buffer_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (dma_buffer_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (dma_buffer_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_dma_buffer_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_dma_buffer_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_dma_buffer_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_dma_buffer_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_dma_buffer_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_dma_buffer_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (dma_buffer_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (dma_buffer_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (dma_buffer_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (dma_buffer_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (dma_buffer_avalon_pixel_source_data)                           //                        .data
	);

	nios_system_dual_clock_fifo dual_clock_fifo (
		.clk_stream_in            (sys_sdram_pll_sys_clk_clk),                                 //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_002_reset_out_reset),                        //         reset_stream_in.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                                   //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_003_reset_out_reset),                        //        reset_stream_out.reset
		.stream_in_ready          (video_alpha_blender_0_avalon_blended_source_ready),         //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_alpha_blender_0_avalon_blended_source_startofpacket), //                        .startofpacket
		.stream_in_endofpacket    (video_alpha_blender_0_avalon_blended_source_endofpacket),   //                        .endofpacket
		.stream_in_valid          (video_alpha_blender_0_avalon_blended_source_valid),         //                        .valid
		.stream_in_data           (video_alpha_blender_0_avalon_blended_source_data),          //                        .data
		.stream_out_ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),             // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket),     //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),       //                        .endofpacket
		.stream_out_valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),             //                        .valid
		.stream_out_data          (dual_clock_fifo_avalon_dc_buffer_source_data)               //                        .data
	);

	nios_system_jtag jtag (
		.clk            (sys_sdram_pll_sys_clk_clk),                            //               clk.clk
		.rst_n          (~rst_controller_004_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	nios_system_nios_custom_instr_floating_point_2_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (processor_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (processor_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (processor_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (processor_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (processor_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (processor_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (processor_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (processor_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (processor_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (processor_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (processor_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (processor_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	nios_system_processor processor (
		.clk                                 (sys_sdram_pll_sys_clk_clk),                               //                       clk.clk
		.reset_n                             (~rst_controller_005_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_005_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (processor_data_master_address),                           //               data_master.address
		.d_byteenable                        (processor_data_master_byteenable),                        //                          .byteenable
		.d_read                              (processor_data_master_read),                              //                          .read
		.d_readdata                          (processor_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (processor_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (processor_data_master_write),                             //                          .write
		.d_writedata                         (processor_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (processor_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (processor_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (processor_instruction_master_address),                    //        instruction_master.address
		.i_read                              (processor_instruction_master_read),                       //                          .read
		.i_readdata                          (processor_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (processor_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (processor_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (processor_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (processor_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_processor_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_processor_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_processor_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_processor_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_processor_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_processor_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_processor_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_processor_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (processor_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (processor_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (processor_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (processor_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (processor_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (processor_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (processor_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (processor_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (processor_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (processor_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (processor_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (processor_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (processor_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (processor_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (processor_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (processor_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (processor_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (processor_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (processor_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (processor_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (processor_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (processor_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (processor_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (processor_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (processor_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (processor_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (processor_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (processor_custom_instruction_master_writerc)              //                          .writerc
	);

	nios_system_rgb_resampler rgb_resampler (
		.clk                      (sys_sdram_pll_sys_clk_clk),                                 //               clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                        //             reset.reset
		.stream_in_startofpacket  (dma_buffer_avalon_pixel_source_startofpacket),              //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (dma_buffer_avalon_pixel_source_endofpacket),                //                  .endofpacket
		.stream_in_valid          (dma_buffer_avalon_pixel_source_valid),                      //                  .valid
		.stream_in_ready          (dma_buffer_avalon_pixel_source_ready),                      //                  .ready
		.stream_in_data           (dma_buffer_avalon_pixel_source_data),                       //                  .data
		.slave_read               (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)                       //                  .data
	);

	nios_system_sdram_controller sdram_controller (
		.clk            (sdram_clk_clk),                                       //   clk.clk
		.reset_n        (~rst_controller_006_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	nios_system_sram_controller sram_controller (
		.clk           (sys_sdram_pll_sys_clk_clk),                                         //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                                //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                           // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                         //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                         //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                         //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                         //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                         //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                         //                   .export
		.address       (mm_interconnect_0_sram_controller_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_controller_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_controller_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_controller_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_controller_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_controller_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_controller_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_system_sys_sdram_pll sys_sdram_pll (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_007_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_sys_clk_clk),          //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_reset_source_reset)    // reset_source.reset
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sys_sdram_pll_sys_clk_clk),                             //           clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_timer_0 timer_0 (
		.clk        (sys_sdram_pll_sys_clk_clk),               //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	nios_system_vga vga (
		.clk           (video_pll_0_vga_clk_clk),                               //                clk.clk
		.reset         (rst_controller_008_reset_out_reset),                    //              reset.reset
		.data          (dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                               // external_interface.export
		.VGA_HS        (vga_HS),                                                //                   .export
		.VGA_VS        (vga_VS),                                                //                   .export
		.VGA_BLANK     (vga_BLANK),                                             //                   .export
		.VGA_SYNC      (vga_SYNC),                                              //                   .export
		.VGA_R         (vga_R),                                                 //                   .export
		.VGA_G         (vga_G),                                                 //                   .export
		.VGA_B         (vga_B)                                                  //                   .export
	);

	nios_system_video_alpha_blender_0 video_alpha_blender_0 (
		.clk                      (sys_sdram_pll_sys_clk_clk),                                          //                    clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                  reset.reset
		.foreground_data          (video_character_buffer_with_dma_0_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),         //                       .ready
		.background_data          (avalon_st_adapter_out_0_data),                                       // avalon_background_sink.data
		.background_startofpacket (avalon_st_adapter_out_0_startofpacket),                              //                       .startofpacket
		.background_endofpacket   (avalon_st_adapter_out_0_endofpacket),                                //                       .endofpacket
		.background_valid         (avalon_st_adapter_out_0_valid),                                      //                       .valid
		.background_ready         (avalon_st_adapter_out_0_ready),                                      //                       .ready
		.output_ready             (video_alpha_blender_0_avalon_blended_source_ready),                  //  avalon_blended_source.ready
		.output_data              (video_alpha_blender_0_avalon_blended_source_data),                   //                       .data
		.output_startofpacket     (video_alpha_blender_0_avalon_blended_source_startofpacket),          //                       .startofpacket
		.output_endofpacket       (video_alpha_blender_0_avalon_blended_source_endofpacket),            //                       .endofpacket
		.output_valid             (video_alpha_blender_0_avalon_blended_source_valid)                   //                       .valid
	);

	nios_system_video_character_buffer_with_dma_0 video_character_buffer_with_dma_0 (
		.clk                  (sys_sdram_pll_sys_clk_clk),                                                                //                       clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                                       //                     reset.reset
		.ctrl_address         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),                               //                          .valid
		.stream_data          (video_character_buffer_with_dma_0_avalon_char_source_data)                                 //                          .data
	);

	nios_system_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_007_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),            //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)      // reset_source.reset
	);

	nios_system_video_scaler video_scaler (
		.clk                      (sys_sdram_pll_sys_clk_clk),                       //                  clk.clk
		.reset                    (rst_controller_001_reset_out_reset),              //                reset.reset
		.stream_in_startofpacket  (rgb_resampler_avalon_rgb_source_startofpacket),   //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_resampler_avalon_rgb_source_endofpacket),     //                     .endofpacket
		.stream_in_valid          (rgb_resampler_avalon_rgb_source_valid),           //                     .valid
		.stream_in_ready          (rgb_resampler_avalon_rgb_source_ready),           //                     .ready
		.stream_in_data           (rgb_resampler_avalon_rgb_source_data),            //                     .data
		.stream_out_ready         (video_scaler_avalon_scaler_source_ready),         // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_avalon_scaler_source_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_avalon_scaler_source_endofpacket),   //                     .endofpacket
		.stream_out_valid         (video_scaler_avalon_scaler_source_valid),         //                     .valid
		.stream_out_data          (video_scaler_avalon_scaler_source_data),          //                     .data
		.stream_out_channel       (video_scaler_avalon_scaler_source_channel)        //                     .channel
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) processor_custom_instruction_master_translator (
		.ci_slave_dataa            (processor_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (processor_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (processor_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (processor_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (processor_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (processor_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (processor_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (processor_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (processor_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (processor_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (processor_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (processor_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (processor_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (processor_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (processor_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (processor_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (processor_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (processor_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (processor_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (processor_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (processor_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (processor_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (processor_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (processor_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (processor_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (processor_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (processor_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (processor_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (processor_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (processor_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (processor_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (processor_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (processor_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (processor_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (processor_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (processor_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (processor_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (processor_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (processor_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (processor_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (processor_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (processor_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (processor_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (processor_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (processor_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (processor_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (processor_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (processor_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (processor_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (processor_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (processor_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (processor_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (processor_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (processor_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (processor_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (processor_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	nios_system_processor_custom_instruction_master_comb_xconnect processor_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (processor_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (processor_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (processor_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (processor_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (processor_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (processor_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (processor_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (processor_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (processor_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (processor_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (processor_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (processor_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (processor_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (processor_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (processor_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (processor_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (processor_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (processor_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (processor_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (processor_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (processor_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (processor_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (processor_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (processor_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) processor_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (processor_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (processor_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (processor_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (processor_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (processor_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (processor_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (processor_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (processor_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (processor_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (processor_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (processor_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (processor_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (processor_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (processor_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (processor_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (processor_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                            // (terminated)
		.ci_master_readrb    (),                                                                            // (terminated)
		.ci_master_writerc   (),                                                                            // (terminated)
		.ci_master_a         (),                                                                            // (terminated)
		.ci_master_b         (),                                                                            // (terminated)
		.ci_master_c         (),                                                                            // (terminated)
		.ci_master_ipending  (),                                                                            // (terminated)
		.ci_master_estatus   (),                                                                            // (terminated)
		.ci_master_clk       (),                                                                            // (terminated)
		.ci_master_clken     (),                                                                            // (terminated)
		.ci_master_reset_req (),                                                                            // (terminated)
		.ci_master_reset     (),                                                                            // (terminated)
		.ci_master_start     (),                                                                            // (terminated)
		.ci_master_done      (1'b0),                                                                        // (terminated)
		.ci_slave_clk        (1'b0),                                                                        // (terminated)
		.ci_slave_clken      (1'b0),                                                                        // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                        // (terminated)
		.ci_slave_reset      (1'b0),                                                                        // (terminated)
		.ci_slave_start      (1'b0),                                                                        // (terminated)
		.ci_slave_done       ()                                                                             // (terminated)
	);

	nios_system_processor_custom_instruction_master_multi_xconnect processor_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (processor_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (processor_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (processor_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (processor_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (processor_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (processor_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (processor_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (processor_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (processor_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (processor_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                         //           .ipending
		.ci_slave_estatus     (),                                                                         //           .estatus
		.ci_slave_clk         (processor_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (processor_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (processor_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (processor_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (processor_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (processor_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (processor_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (processor_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (processor_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (processor_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (processor_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (processor_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (processor_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (processor_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (processor_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (processor_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (processor_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (processor_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (processor_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (processor_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (processor_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (processor_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (processor_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (processor_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) processor_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (processor_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (processor_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (processor_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (processor_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (processor_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (processor_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (processor_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (processor_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (processor_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (processor_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (processor_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (processor_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (processor_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (processor_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (processor_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (processor_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (processor_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (processor_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (processor_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (processor_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (processor_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (processor_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (processor_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (processor_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (processor_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (processor_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                                // (terminated)
		.ci_master_readrb    (),                                                                                // (terminated)
		.ci_master_writerc   (),                                                                                // (terminated)
		.ci_master_a         (),                                                                                // (terminated)
		.ci_master_b         (),                                                                                // (terminated)
		.ci_master_c         (),                                                                                // (terminated)
		.ci_master_ipending  (),                                                                                // (terminated)
		.ci_master_estatus   ()                                                                                 // (terminated)
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_sdram_clk_clk                                            (sdram_clk_clk),                                                                            //                                     sys_sdram_pll_sdram_clk.clk
		.sys_sdram_pll_sys_clk_clk                                              (sys_sdram_pll_sys_clk_clk),                                                                //                                       sys_sdram_pll_sys_clk.clk
		.dma_buffer_reset_reset_bridge_in_reset_reset                           (rst_controller_001_reset_out_reset),                                                       //                      dma_buffer_reset_reset_bridge_in_reset.reset
		.jtag_reset_reset_bridge_in_reset_reset                                 (rst_controller_004_reset_out_reset),                                                       //                            jtag_reset_reset_bridge_in_reset.reset
		.processor_reset_reset_bridge_in_reset_reset                            (rst_controller_005_reset_out_reset),                                                       //                       processor_reset_reset_bridge_in_reset.reset
		.sdram_controller_reset_reset_bridge_in_reset_reset                     (rst_controller_006_reset_out_reset),                                                       //                sdram_controller_reset_reset_bridge_in_reset.reset
		.dma_buffer_avalon_pixel_dma_master_address                             (dma_buffer_avalon_pixel_dma_master_address),                                               //                          dma_buffer_avalon_pixel_dma_master.address
		.dma_buffer_avalon_pixel_dma_master_waitrequest                         (dma_buffer_avalon_pixel_dma_master_waitrequest),                                           //                                                            .waitrequest
		.dma_buffer_avalon_pixel_dma_master_read                                (dma_buffer_avalon_pixel_dma_master_read),                                                  //                                                            .read
		.dma_buffer_avalon_pixel_dma_master_readdata                            (dma_buffer_avalon_pixel_dma_master_readdata),                                              //                                                            .readdata
		.dma_buffer_avalon_pixel_dma_master_readdatavalid                       (dma_buffer_avalon_pixel_dma_master_readdatavalid),                                         //                                                            .readdatavalid
		.dma_buffer_avalon_pixel_dma_master_lock                                (dma_buffer_avalon_pixel_dma_master_lock),                                                  //                                                            .lock
		.processor_data_master_address                                          (processor_data_master_address),                                                            //                                       processor_data_master.address
		.processor_data_master_waitrequest                                      (processor_data_master_waitrequest),                                                        //                                                            .waitrequest
		.processor_data_master_byteenable                                       (processor_data_master_byteenable),                                                         //                                                            .byteenable
		.processor_data_master_read                                             (processor_data_master_read),                                                               //                                                            .read
		.processor_data_master_readdata                                         (processor_data_master_readdata),                                                           //                                                            .readdata
		.processor_data_master_readdatavalid                                    (processor_data_master_readdatavalid),                                                      //                                                            .readdatavalid
		.processor_data_master_write                                            (processor_data_master_write),                                                              //                                                            .write
		.processor_data_master_writedata                                        (processor_data_master_writedata),                                                          //                                                            .writedata
		.processor_data_master_debugaccess                                      (processor_data_master_debugaccess),                                                        //                                                            .debugaccess
		.processor_instruction_master_address                                   (processor_instruction_master_address),                                                     //                                processor_instruction_master.address
		.processor_instruction_master_waitrequest                               (processor_instruction_master_waitrequest),                                                 //                                                            .waitrequest
		.processor_instruction_master_read                                      (processor_instruction_master_read),                                                        //                                                            .read
		.processor_instruction_master_readdata                                  (processor_instruction_master_readdata),                                                    //                                                            .readdata
		.processor_instruction_master_readdatavalid                             (processor_instruction_master_readdatavalid),                                               //                                                            .readdatavalid
		.dma_buffer_avalon_control_slave_address                                (mm_interconnect_0_dma_buffer_avalon_control_slave_address),                                //                             dma_buffer_avalon_control_slave.address
		.dma_buffer_avalon_control_slave_write                                  (mm_interconnect_0_dma_buffer_avalon_control_slave_write),                                  //                                                            .write
		.dma_buffer_avalon_control_slave_read                                   (mm_interconnect_0_dma_buffer_avalon_control_slave_read),                                   //                                                            .read
		.dma_buffer_avalon_control_slave_readdata                               (mm_interconnect_0_dma_buffer_avalon_control_slave_readdata),                               //                                                            .readdata
		.dma_buffer_avalon_control_slave_writedata                              (mm_interconnect_0_dma_buffer_avalon_control_slave_writedata),                              //                                                            .writedata
		.dma_buffer_avalon_control_slave_byteenable                             (mm_interconnect_0_dma_buffer_avalon_control_slave_byteenable),                             //                                                            .byteenable
		.jtag_avalon_jtag_slave_address                                         (mm_interconnect_0_jtag_avalon_jtag_slave_address),                                         //                                      jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                                           (mm_interconnect_0_jtag_avalon_jtag_slave_write),                                           //                                                            .write
		.jtag_avalon_jtag_slave_read                                            (mm_interconnect_0_jtag_avalon_jtag_slave_read),                                            //                                                            .read
		.jtag_avalon_jtag_slave_readdata                                        (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                                        //                                                            .readdata
		.jtag_avalon_jtag_slave_writedata                                       (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                                       //                                                            .writedata
		.jtag_avalon_jtag_slave_waitrequest                                     (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),                                     //                                                            .waitrequest
		.jtag_avalon_jtag_slave_chipselect                                      (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                                      //                                                            .chipselect
		.processor_debug_mem_slave_address                                      (mm_interconnect_0_processor_debug_mem_slave_address),                                      //                                   processor_debug_mem_slave.address
		.processor_debug_mem_slave_write                                        (mm_interconnect_0_processor_debug_mem_slave_write),                                        //                                                            .write
		.processor_debug_mem_slave_read                                         (mm_interconnect_0_processor_debug_mem_slave_read),                                         //                                                            .read
		.processor_debug_mem_slave_readdata                                     (mm_interconnect_0_processor_debug_mem_slave_readdata),                                     //                                                            .readdata
		.processor_debug_mem_slave_writedata                                    (mm_interconnect_0_processor_debug_mem_slave_writedata),                                    //                                                            .writedata
		.processor_debug_mem_slave_byteenable                                   (mm_interconnect_0_processor_debug_mem_slave_byteenable),                                   //                                                            .byteenable
		.processor_debug_mem_slave_waitrequest                                  (mm_interconnect_0_processor_debug_mem_slave_waitrequest),                                  //                                                            .waitrequest
		.processor_debug_mem_slave_debugaccess                                  (mm_interconnect_0_processor_debug_mem_slave_debugaccess),                                  //                                                            .debugaccess
		.rgb_resampler_avalon_rgb_slave_read                                    (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_read),                                    //                              rgb_resampler_avalon_rgb_slave.read
		.rgb_resampler_avalon_rgb_slave_readdata                                (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_readdata),                                //                                                            .readdata
		.sdram_controller_s1_address                                            (mm_interconnect_0_sdram_controller_s1_address),                                            //                                         sdram_controller_s1.address
		.sdram_controller_s1_write                                              (mm_interconnect_0_sdram_controller_s1_write),                                              //                                                            .write
		.sdram_controller_s1_read                                               (mm_interconnect_0_sdram_controller_s1_read),                                               //                                                            .read
		.sdram_controller_s1_readdata                                           (mm_interconnect_0_sdram_controller_s1_readdata),                                           //                                                            .readdata
		.sdram_controller_s1_writedata                                          (mm_interconnect_0_sdram_controller_s1_writedata),                                          //                                                            .writedata
		.sdram_controller_s1_byteenable                                         (mm_interconnect_0_sdram_controller_s1_byteenable),                                         //                                                            .byteenable
		.sdram_controller_s1_readdatavalid                                      (mm_interconnect_0_sdram_controller_s1_readdatavalid),                                      //                                                            .readdatavalid
		.sdram_controller_s1_waitrequest                                        (mm_interconnect_0_sdram_controller_s1_waitrequest),                                        //                                                            .waitrequest
		.sdram_controller_s1_chipselect                                         (mm_interconnect_0_sdram_controller_s1_chipselect),                                         //                                                            .chipselect
		.sram_controller_avalon_sram_slave_address                              (mm_interconnect_0_sram_controller_avalon_sram_slave_address),                              //                           sram_controller_avalon_sram_slave.address
		.sram_controller_avalon_sram_slave_write                                (mm_interconnect_0_sram_controller_avalon_sram_slave_write),                                //                                                            .write
		.sram_controller_avalon_sram_slave_read                                 (mm_interconnect_0_sram_controller_avalon_sram_slave_read),                                 //                                                            .read
		.sram_controller_avalon_sram_slave_readdata                             (mm_interconnect_0_sram_controller_avalon_sram_slave_readdata),                             //                                                            .readdata
		.sram_controller_avalon_sram_slave_writedata                            (mm_interconnect_0_sram_controller_avalon_sram_slave_writedata),                            //                                                            .writedata
		.sram_controller_avalon_sram_slave_byteenable                           (mm_interconnect_0_sram_controller_avalon_sram_slave_byteenable),                           //                                                            .byteenable
		.sram_controller_avalon_sram_slave_readdatavalid                        (mm_interconnect_0_sram_controller_avalon_sram_slave_readdatavalid),                        //                                                            .readdatavalid
		.sysid_qsys_0_control_slave_address                                     (mm_interconnect_0_sysid_qsys_0_control_slave_address),                                     //                                  sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                    (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                                    //                                                            .readdata
		.timer_0_s1_address                                                     (mm_interconnect_0_timer_0_s1_address),                                                     //                                                  timer_0_s1.address
		.timer_0_s1_write                                                       (mm_interconnect_0_timer_0_s1_write),                                                       //                                                            .write
		.timer_0_s1_readdata                                                    (mm_interconnect_0_timer_0_s1_readdata),                                                    //                                                            .readdata
		.timer_0_s1_writedata                                                   (mm_interconnect_0_timer_0_s1_writedata),                                                   //                                                            .writedata
		.timer_0_s1_chipselect                                                  (mm_interconnect_0_timer_0_s1_chipselect),                                                  //                                                            .chipselect
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //  video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                                                            .write
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                                                            .read
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                                                            .readdata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                                                            .writedata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //                                                            .byteenable
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                                                            .waitrequest
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                                                            .chipselect
		.video_character_buffer_with_dma_0_avalon_char_control_slave_address    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // video_character_buffer_with_dma_0_avalon_char_control_slave.address
		.video_character_buffer_with_dma_0_avalon_char_control_slave_write      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                                                            .write
		.video_character_buffer_with_dma_0_avalon_char_control_slave_read       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                                                            .read
		.video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                                                            .readdata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                                                            .writedata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                                                            .byteenable
		.video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect)  //                                                            .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_sys_clk_clk),          //       clk.clk
		.reset         (rst_controller_005_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (processor_irq_irq)                   //    sender.irq
	);

	nios_system_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (2),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sys_sdram_pll_sys_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),              // in_rst_0.reset
		.in_0_data           (video_scaler_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (video_scaler_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (video_scaler_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (video_scaler_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (video_scaler_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (video_scaler_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                    //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                   //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                   //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),           //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)              //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                   // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset), // reset_in1.reset
		.clk            (),                                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset),   // reset_in1.reset
		.clk            (sys_sdram_pll_sys_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (sys_sdram_pll_sys_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset),   // reset_in1.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (rst_controller_reset_out_reset),     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (sys_sdram_pll_reset_source_reset),   // reset_in2.reset
		.clk            (sys_sdram_pll_sys_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (processor_debug_reset_request_reset),    // reset_in1.reset
		.reset_in2      (sys_sdram_pll_reset_source_reset),       // reset_in2.reset
		.clk            (sys_sdram_pll_sys_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_005_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset),   // reset_in1.reset
		.clk            (sdram_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset),   // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (rst_controller_reset_out_reset),     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (sys_sdram_pll_reset_source_reset),   // reset_in2.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
